library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
use UNISIM.vcomponents.all;


entity attitude_calc is
	port (
		clk : in  STD_LOGIC;
		read_regs : in  STD_LOGIC_VECTOR (143 downto 0);
		write_en : out  STD_LOGIC;
		write_addr : out  STD_LOGIC_VECTOR (7 downto 0);
		write_data : out  STD_LOGIC_VECTOR (15 downto 0)
	);
end attitude_calc;

architecture Behavioral of attitude_calc is
	constant ax_offset: std_logic_vector(17 downto 0) := signed(-430);
	constant ay_offset: std_logic_vector(17 downto 0) := signed(8);
	constant az_offset: std_logic_vector(17 downto 0) := signed(85);
	
	constant gx_offset: std_logic_vector(17 downto 0) := signed(32);
	constant gy_offset: std_logic_vector(17 downto 0) := signed(28);
	constant gz_offset: std_logic_vector(17 downto 0) := signed(4);


	constant Dt: std_logic_vector(17 downto 0) := "010100011110101110"; -- * 2^-25 = 0.0025; Time constant in s
	constant Kd: std_logic_vector(17 downto 0) := "011111001110000011"; --0.9756098, 1 integer place; depends on Dt
	constant Kp: std_logic_vector(17 downto 0) := "000000110001111101"; --0.0243902, 1 integer place depends on Dt
	
	--Scale gyro readings from 65.5 lsb/(deg/s) to milliradians/s
	--TODO: change gyro range on uProc to +-500deg
	--Also increase sampling rate, forsrs
	constant gyro_scale: std_logic_vector(17 downto 0) := "010001000011011011"-- * 2^-18 = 0.266462;
	

	signal ax_raw, ayraw, azraw: std_logic_vector(17 downto 0);
	signal axc, ayc, azc: std_logic_vector(17 downto 0);
	signal acc_pitch, acc_roll: std_logic_vector(17 downto 0);
		
	signal gx_raw, gy_raw, gz_raw: std_logic_vector(17 downto 0); --*2^0
	signal gx, gy, gz: std_logic_vector(17 downto 0); --todo: find exponent for this
	signal gx_int, gy_int: std_logic_vector(17 downto 0);
	
	
	signal last_pitch, last_roll: std_logic_vector(17 downto 0);
	signal p_pitch, d_pitch: std_logic_vector(17 downto 0);	
	signal p_roll, d_roll: std_logic_vector(17 downto 0);
	signal pitch, roll: std_logic_vector(17 downto 0);
	signal m_pitch, m_roll: std_logic_vector(17 downto 0);

	signal atan_rdy1, atan_rdy2: std_logic;
	
	
	component arctan
		port (
			x_in : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			y_in : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			phase_out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			rdy : OUT STD_LOGIC;
			clk : IN STD_LOGIC
		);
	end component;

begin

	--=======================--
	-- Load data from register file (and sign-extend)
	ax_raw <= std_logic_vector(resize(signed(read_regs(15 downto 0)), 18));
	ay_raw <= std_logic_vector(resize(signed(read_regs(31 downto 16)), 18));
	az_raw <= std_logic_vector(resize(signed(read_regs(47 downto 32)), 18));
	
	gx_raw <= std_logic_vector(resize(signed(read_regs(63 downto 48)), 18));
	gy_raw <= std_logic_vector(resize(signed(read_regs(79 downto 64)), 18));
	gz_raw <= std_logic_vector(resize(signed(read_regs(95 downto 80)), 18));
	
	
	--=======================--
	-- Gyro processing section
	-- Pitch:
	
	--Preadd-multiply: op=0x11; P=a*(b+d) = (gx_raw + gx_offset) * gx_scale
	dsp_gx1: entity work.dsp48a1_wrapper(Behavioral)
		port map(
			a => gyro_scale,
			b => gx_raw,
			d => gx_offset,
			p => gx,
			
			rst => rst,
			clk => clk,
			clk_en => clk_en,
			opmode => X"11"	
		);
	
	--Multiply-postadd: op=0x1D; P=c+(a*b) = (gx * Dt) + last_pitch
	dsp_gx2: entity work.dsp48a1_wrapper(Behavioral)
		port map(
			a => gx(,
			b => Dt,
			c => last_pitch,
			p => gx_int,
			
			rst => rst,
			clk => clk,
			clk_en => clk_en,
			opmode => X"1D"	
		);
		
	--Multiply: op=0x01; C_P_out=a*b = gx_int * Kp (cascade to dsp_pitch)
	dsp_p_pitch: entity work.dsp48a1_wrapper(Behavioral)
		port map(
			a => gx_int,
			b => Kp,
			c_p_out => p_pitch,
			
			rst => rst,
			clk => clk,
			clk_en => clk_en,
			opmode => X"01"	
		);
		
		
	------------------------
	--Roll:

	--Preadd-multiply: op=0x11; P=a*(b+d) = (gy_raw + gy_offset) * gy_scale
	dsp_gy1: entity work.dsp48a1_wrapper(Behavioral)
		port map(
			a => gyro_scale,
			b => gy_raw,
			d => gy_offset,
			p => gy,
			
			rst => rst,
			clk => clk,
			clk_en => clk_en,
			opmode => X"11"
		);
	
	--Multiply-postadd: op=0x1D; P=c+(a*b) = (gy * Dt) + last_roll
	dsp_gy2: entity work.dsp48a1_wrapper(Behavioral)
		port map(
			a => gy,
			b => Dt,
			c => last_roll,
			p => gy_int,
			
			rst => rst,
			clk => clk,
			clk_en => clk_en,
			opmode => X"1D"	
		);
	
	--Multiply: op=0x01; C_P_out=a*b = gy_int * Kp (cascade to dsp_roll)
	dsp_p_roll: entity work.dsp48a1_wrapper(Behavioral)
		port map(
			a => gy_int,
			b => Kp,
			c_p_out => p_roll,
			
			rst => rst,
			clk => clk,
			clk_en => clk_en,
			opmode => X"01"	
		);
	
	
	
	--=========================--
	-- Accelerometer section
	
	--Add stage: add constants to raw sensor values
	axc <= signed(ax_raw) + signed(ax_offset);
	ayc <= signed(ay_raw) + signed(ay_offset);
	azc <= signed(az_raw) + signed(az_offset);
	
	--Trig stage: take arctangent of offset sensor values
	arctan_i1: arctan
		port map(
			x_in => axc,
			y_in => azc,
			phase_out => acc_pitch,
			rdy => atan_rdy1,
			clk => clk
		);
		
	arctan_i2: arctan
		port map(
			x_in => ayc,
			y_in => azc,
			phase_out => acc_roll,
			rdy => atan_rdy2,
			clk => clk
		);
	
	
	
	
	--=========================--
	-- Combine gyro and accelerometer data
	
	--Cascade multiply-postadd: op=0x05; P=P_in+(a*b) = (atan_out1 * Kd) + p_pitch
	dsp_pitch: entity work.dsp48a1_wrapper(Behavioral)
		port map(
			a => acc_pitch,
			b => Kd,
			c_p_in => p_pitch,
			p => pitch,
			
			rst => rst,
			clk => clk,
			clk_en => clk_en,
			opmode => X"05"	
		);
		
	--Cascade multiply-postadd: op=0x05; P=P_in+(a*b) = (atan_out2 * Kd) + p_roll
	dsp_roll: entity work.dsp48a1_wrapper(Behavioral)
		port map(
			a => acc_roll,
			b => Kd,
			c_p_in => p_roll,
			p => roll,
			
			rst => rst,
			clk => clk,
			clk_en => clk_en,
			opmode => X"05"	
		);
	
	--Add stage: correct for mounting angle
	m_pitch <= signed(pitch) + signed(pitch_corr);
	m_roll <= signed(roll) + signed(roll_corr);
	
	





end Behavioral;

